/*******************************************************************
* Module Name: SPI Flash controller
* 
* Description: 
* This module [briefly describe the module's purpose and functionality].
* [Optional: Additional notes on functionality, special cases, or constraints.]
*
* Inputs:
* clk - 1-bit clock input signal for synchronizing the module's operations.
* rstn - 1-bit active low reset signal for initializing or resetting the module's internal state.
* [Document other inputs here if applicable...]
*
* Outputs:
* [Document outputs here if applicable...]
*
* Author: Tin Sorić
* Date: [Date, e.g., "YYYY-MM-DD"]
*******************************************************************/


module spi_flash (
    input   clk,
    input   rstn
);


endmodule